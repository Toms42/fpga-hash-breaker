module pad_tester